//top test